CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 108 189 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7876 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 1023 203 0 18 19
10 8 7 6 5 4 3 2 18 19
1 1 1 0 0 1 1 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
6369 0 0
2
43530.4 1
0
9 2-In AND~
219 540 53 0 3 22
0 14 10 13
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9172 0 0
2
43530.4 2
0
9 2-In AND~
219 390 52 0 3 22
0 12 11 14
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7100 0 0
2
43530.4 3
0
6 74112~
219 604 225 0 7 32
0 17 13 15 13 17 20 9
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3820 0 0
2
43530.4 4
0
6 74112~
219 504 226 0 7 32
0 17 14 15 14 17 21 10
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
7678 0 0
2
43530.4 5
0
6 74112~
219 395 231 0 7 32
0 17 12 15 12 17 22 11
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
961 0 0
2
43530.4 6
0
6 74112~
219 289 231 0 7 32
0 17 16 15 16 17 23 12
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3178 0 0
2
43530.4 7
0
6 74LS48
188 848 235 0 14 29
0 9 10 11 12 24 25 2 3 4
5 6 7 8 26
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
43530.4 8
0
2 +V
167 131 125 0 1 3
0 17
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
43530.4 9
0
7 Pulser~
4 70 313 0 10 12
0 27 28 15 29 0 0 5 5 4
7
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8885 0 0
2
43530.4 10
0
38
7 7 2 0 0 4224 0 9 2 0 0 5
880 199
973 199
973 272
1038 272
1038 239
8 6 3 0 0 4224 0 9 2 0 0 5
880 208
978 208
978 267
1032 267
1032 239
9 5 4 0 0 4224 0 9 2 0 0 5
880 217
983 217
983 262
1026 262
1026 239
10 4 5 0 0 4224 0 9 2 0 0 5
880 226
988 226
988 257
1020 257
1020 239
11 3 6 0 0 4224 0 9 2 0 0 5
880 235
993 235
993 247
1014 247
1014 239
12 2 7 0 0 4224 0 9 2 0 0 3
880 244
1008 244
1008 239
13 1 8 0 0 4224 0 9 2 0 0 3
880 253
1002 253
1002 239
7 1 9 0 0 4224 0 5 9 0 0 4
628 189
803 189
803 199
816 199
0 2 10 0 0 12416 0 0 9 14 0 6
539 184
560 184
560 247
798 247
798 208
816 208
0 3 11 0 0 4224 0 0 9 18 0 4
433 243
803 243
803 217
816 217
0 4 12 0 0 4224 0 0 9 26 0 4
327 155
808 155
808 226
816 226
0 4 13 0 0 4096 0 0 5 13 0 3
566 95
566 207
580 207
3 2 13 0 0 8320 0 3 5 0 0 4
561 53
566 53
566 189
580 189
2 7 10 0 0 0 0 3 6 0 0 6
516 62
512 62
512 159
539 159
539 190
528 190
0 4 14 0 0 4224 0 0 6 17 0 3
429 52
429 208
480 208
0 1 14 0 0 0 0 0 3 17 0 3
465 52
465 44
516 44
3 2 14 0 0 0 0 4 6 0 0 4
411 52
466 52
466 190
480 190
2 7 11 0 0 0 0 4 7 0 0 6
366 61
356 61
356 248
433 248
433 195
419 195
1 0 12 0 0 0 0 4 0 0 25 3
366 43
335 43
335 195
3 0 15 0 0 8192 0 5 0 0 23 3
574 198
570 198
570 304
3 0 15 0 0 0 0 6 0 0 23 3
474 199
470 199
470 304
3 0 15 0 0 0 0 7 0 0 23 3
365 204
361 204
361 304
0 0 15 0 0 4224 0 0 0 27 0 2
251 304
690 304
0 4 12 0 0 0 0 0 7 25 0 3
343 195
343 213
371 213
0 2 12 0 0 0 0 0 7 26 0 2
326 195
371 195
7 0 12 0 0 0 0 8 0 0 0 3
313 195
327 195
327 94
3 3 15 0 0 0 0 11 8 0 0 4
94 304
251 304
251 204
259 204
0 4 16 0 0 8192 0 0 8 29 0 3
144 189
144 213
265 213
1 2 16 0 0 4224 0 1 8 0 0 4
120 189
251 189
251 195
265 195
5 0 17 0 0 4096 0 8 0 0 38 2
289 243
289 274
5 0 17 0 0 4096 0 5 0 0 38 2
604 237
604 274
5 0 17 0 0 0 0 6 0 0 38 2
504 238
504 274
5 0 17 0 0 0 0 7 0 0 38 2
395 243
395 274
0 1 17 0 0 0 0 0 5 38 0 2
604 134
604 162
0 1 17 0 0 0 0 0 6 38 0 2
504 134
504 163
1 0 17 0 0 0 0 7 0 0 38 2
395 168
395 134
0 1 17 0 0 0 0 0 8 38 0 3
287 134
289 134
289 168
1 0 17 0 0 4224 0 10 0 0 0 4
131 134
691 134
691 274
131 274
1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
239 359 396 383
249 367 385 383
17 AMOLATO, JENEVEVE
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
